tree decoder